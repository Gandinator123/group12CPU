module mips_cpu_harvard();
logic a;

logic b;
endmodule