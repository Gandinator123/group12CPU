module mips_cpu_harvard();


endmodule