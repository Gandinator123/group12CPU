module mips_cpu_harvard();

input a;
endmodule