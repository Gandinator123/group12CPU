module mips_cpu_harvard();
logic a;

logic b;

logic c;

logic d;

endmodule