module mips_cpu_harvard();
logic a;

endmodule