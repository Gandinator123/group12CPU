module mips_cpu_harvard();
logic a;

logic b;

logic ccc;

logic rohan;
logic d;


endmodule